


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity datapath is
	port(
		CLK, RST: in std_logic;
			-- data inputs
			-- data outputs
			-- control signals
			-- status signals
		);
entity datapath;